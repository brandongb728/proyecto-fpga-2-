LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL; 

ENTITY Display IS 
PORT (
	numero   : IN INTEGER RANGE 0 TO 9;
	SEG7 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)  
);
END ENTITY;
 
ARCHITECTURE behaviour OF Display IS
BEGIN
display_output : PROCESS(numero)
BEGIN
	CASE numero IS
	 WHEN 0 =>
		SEG7 <= B"1000000";
	 WHEN 1 =>
		SEG7 <= B"1111001";
	 WHEN 2 =>
		SEG7 <= B"0100100";
	 WHEN 3 =>
		SEG7 <= B"0110000";
	 WHEN 4 =>
		SEG7 <= B"0011001";
	 WHEN 5 =>
		SEG7 <= B"0010010";
	 WHEN 6 =>
		SEG7 <= B"0000010";
	 WHEN 7 =>
		SEG7 <= B"1111000";
	 WHEN 8 =>
		SEG7 <= B"0000000";
	 WHEN 9 =>
		SEG7 <= B"0010000";
	 WHEN OTHERS =>
		SEG7 <= B"0000000"; 
	END CASE; 	
END PROCESS;
END ARCHITECTURE;